module bool_tb();
